module None();

endmodule