module Wall();
endmodule