module Seven_Segment(i, a, b, c, d, e, f, g);
	input [3:0]i;
	output a, b, c, d, e, f, g;
	
assign a = ~((i[0] & ~i[1] & ~i[2]) | (i[0] & ~i[3]) | (i[1] & i[2]) | (~i[0] & i[2]) | (~i[0] & ~i[1] & ~i[3]) | (~i[0] & i[1] & i[3]));
assign b = ~((~i[0] & ~i[1]) | (~i[1] & ~i[3]) | (i[0] & ~i[2] & i[3]) | (~i[0] & ~i[2] & ~i[3]) | (~i[0] & i[2] & i[3]));
assign c = ~((~i[0] & i[3]) | (~i[0] & ~i[2]) | (~i[2] & i[3]) | (i[0] & ~i[1]) | (i[1] & ~i[0]));
assign d = ~((i[0] & ~i[2]) | (i[1] & ~i[2] & i[3]) | (~i[0] & ~i[1] & ~i[3]) | (i[1] & i[2] & ~i[3]) | (~i[1] & i[2] & i[3]));
assign e = ~((~i[1] & ~i[3]) | (i[0] & i[1]) | (i[0] & i[2]) | (i[2] & ~i[3]));
assign f = ~((~i[2] & ~i[3]) | (~i[0] & i[1] & ~i[2]) | (i[1] & ~i[3]) | (i[0] & ~i[1]) | (i[0] & i[2]));
assign g = ~((~i[0] & i[1] & ~i[2]) | (i[0] & i[3]) | (i[0] & ~i[1]) | (i[2] & ~i[3]) | (~i[1] & i[2]));	

endmodule
