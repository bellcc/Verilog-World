module Wall(color);
endmodule