module Blank();

endmodule