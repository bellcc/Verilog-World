module Blank(in, out);

input in;
output out;

endmodule
