module Scooter(color);
endmodule