module myModule(in, out);
	input in;
	output out;
	
	//Test myTest(in, in, out);
	
	assign out = in;
endmodule