module Blank(in, out);
endmodule