module Wall(color);
	output [23:0]color;
	
	assign color = 24'hFF0000;
endmodule